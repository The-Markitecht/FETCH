
        `timescale 1 ns / 1 ns

        module visor_program (
            clock_ifc clk,
            code_ifc code
        );
            assign code.content = 
    
